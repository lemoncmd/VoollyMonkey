module main

import ast
import token

fn main() {
}
